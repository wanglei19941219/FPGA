module sdram_wr_module(
        input                   s_clk                   ;
        input                   s_rst_n                 ;
                                                                                                                                                                                                                       


);





































endmodule
