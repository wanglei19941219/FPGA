// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
hEUpJa/6oe1pvxMHtBhinFCt4CjW3lGsd9kHHAUfnUNuoGv4yEbRCDg/SROvJ46D0nfagtiDPKux
ZBUTKqm+4oK76WgVzMxXaCHL3yG2OiPmWqwCsKcZei6+jAM8mMn5uhv3KQp9IU2qM3JL2h+pt2/P
XsHrJldtxOdG6skyUYT964nb4lxLCOKAR3RvPUVDoqAmWe66kF5tSjuuiGHkHTRInWPf04pT3EwL
M1ufnTFTkVTqXWsQyJ3a2qT++ThefQ7E7p8itIe9sWZBcyYuLcU962CbgsDjcG+4n37TbmCogEU0
PjN4JPDuhom1PM5e2dXj/JJ4Qw29lAUwIzMZLA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
TBhwoJcV/NInaGqe0HegbGQL1AW/ilNxfUQv/Z82NO6tm7OcY3nVk4E1/yKucCPKbFn85tB6MecO
TmgUvE575X0fJcffIhl7g0/BOM74IQHb5n4mlHIpDVun+H+h6M99qNoe7Pk+EttFQBDJZMLWuB9o
2vnsPiDZ+mcAu+TAWpKA4fOV5FxBcA09XXNGy5KL9xIeh4ZGU4JSmMmcnbDTucC51XAvtaRsaDhV
mS6LmeFgku7jM6Jw9BnjoMppBPnWrLY4ODymH5YX9fqe0y0ieCraoRchNYP1OajwYg80DapkgAcz
k6wCZYFJoFgX6LD/92N4anUthqYxPlH2UxqqzllZHQKnraAvXMbBp+S6+cdVWDUZAzcjFWnNZxVV
FMgmj6lQCd8C/zS6Q7RVYl312nUDhiiJGUJAI61nQHrWuyvlX6gaQGQi2ItuZnHw2U72rYVDxtWY
uKsDEGObzsMeK6yeixT5PX10L392DuAuuZWPoroGblprIMbJHgpPF0HpFiPQNJNMhoVOgYSi8upi
vXGCGajPRsGb4iEnECwNLTu2MvE4EyZX8uJKSL7I/e/gxkVf8YceY+PouLMQRrQ5Lh5kHRjoHkgc
vQNsnaTLZ7G48uv6Bm/FtnAAeL3pA/Dcwi2OaawHmDrQwinzhMhufIGsQ5aD4S6TSkUi1+GC0079
V/rYf6azEdxbs1ILi8eZKveVumMqOmRQ651v/PDW+EGFELCRFsXl+g7FUJ16ro/kii8dK0w9yjIX
D7Iqf6LHq3+ef5J5eOo+b9pD5AIEItOXb74d9aBlCiMxrTF05pt0wiVp/uXwW9Cv9EuziNS/5kFu
FXfacuKZZs5H7Zunzo5BLemkjf6nSPO0lC5yarrYUHN5UcezIcC4XyB+aExAGptaQeBJfO2p7YQJ
IeA5grmSaqsEob2vrtkIUqS1hWCo5Dc/rNjknlFkF/zNHbyK7XPJIK8SYgRanOiHSkCW+efi2rGv
d96d4dgD6E7eNq5ax8BIbOFRytglQIEWXDYHv22g9KS0rDmlfmNbxXeol4/xUoOXr4uxkA0wLCbO
SQ+4MrH+gpyWTJeFKCoBPHHSFrkqO/200Zd2rhFJi1kaUpY55ntN2y+QLz0ZyibR+PXDvbVITlbh
O7mKqqqa+EHBEZt2ng/CWh3pFrDexILXC/44txVDJQT3VmAT0f0wStchbL776QuiQKPOjReCaaQp
Cd5Q+h/OcItSzyc2vPtxzxo1T2yIjTwT1Fzq1kx4K/0ueTPB0r/3rGMVKpGEX9EJlkpNDV6e+I4O
PesVpd64eNzAiqwKAC5dCL7LYAfnXgIdtAQ2MUidFZonRYcvS2jQL+5q2Erz0mtu19BYe8x9qiOs
YFHQnjAXjHh/xVa2n7lBxLLSIDnzfcG/lk+Lm1gPNSVfw8E7mn/b8R2EkwLE2euKggZQkRjzMviY
lkVvmoPCc50boZX24K9xRNjAoLzhq14Of9sSEJJN15BBlI2eJBu2Gui4V0gvpcwOWrHvYjp9EB3l
ESseWHOEgFsA/xJzutnd3TYxyvP1ZvF28CxgGAydSuoD4gSTRhldlYN468oR/axantZw51nK+f8z
vM6TtnCw2/N3em30/e2yOd4t78fsYczlja0G3ZqKLwMI81JeGybOiWgKrAAOjSFwY94/MAkDE99w
cLzHIfmyU10h7vedrRa9i48gJWBIvlM2sTViM5ATM3lsC/V3kyZqVOAQc7XBSqSdF1QfqbSspI6i
DKi1UYU9KkRH8HOdaWgSzFUvlY+jwt9YYP9FIIOkiGxuYN6EnH9e4S5x4uP4nmns2492s6E7BSIO
m9efcr5b8c7K7j+aOD2YLdsOH3sUd9+o/Nm9v9XdLDxco6CMCZljZv/vPW5mq4ztMUWRnc1vCXdf
3nt4/HHaVUTjXmVR3FCyetq587uB/UTECJ5FBcINmYYHnNxbJyiZ72v/W3SeRYvPaHeUJlmbyEJu
+NLzLEeT76pNDriHT8znODKV6DQ+Bbz9rjj5zTxCRVIuIvc8F/lOUluxa3Uktzn+9WKop/c7H2q/
NlmfD5r+bteHYxyLgb5OCSEQCko7Knfeu52HaHVEvK0WBL7jc+FRXQLyhaouYyypqrFz8cZsNn02
pIhoT4GB6AF3MdkK0OJ6Mj4+3B3l+86P8bE1hedgWhgeP/VdRWOONtlkKhBZ0b/vwwxZq+jV2AfR
8kPJa+K3xTj2usHmiiqo1OL9GrYlc+2LAkP6g0IQ1/bYR2HgFMSC/SdR9f8/8fd407P77y95aikk
A2G7cf/q7K1V2VsR3g1rvcnBO6i/UBpAcwIY20UN3Rr2NatsFEGYKy3onjgrpJMMT9Bcrn/F7UtN
UTeKIaYTovhWcLgcBVLEp6/+OFyQpgwKx6H19/yQkyylR623BRYLtc8PzPbEu+T1t5JFJVyy0mdN
9t0wuEmkfvA/O4hmCrYcVJGDEYqN5Cjj3YEcuFVo+CkW3QFhyQjqVkb9DwnqR9O/LW5IV+MhusmH
SD5XSnRaYZdvCXsQ5oRRFvJPDSHa0rxvBT5AhbPkyUfkdcbjEOIJALqAECIbE8q4AtDmaz3hjpZg
waXIAogmCnIMldUgz3K9gKhhPSd4ueTg2Qea4jUWug54bXQPmnk1dNZD9jUlHEWnT8AWsEiAInQl
iNP6UR73TLU6HmDtJ0Ng2PW0YLtUKE0EyHkpWpCwY+EDL6CSgASGdnUiv0rhQKjhTBfi+7HjRXuv
oNUErmhW5HZrv542DymN1kn7eQ1qSVixzMpokspUtB5g1ZKM4eiRz+LaV5kBPpRbIypFd2K+kpS5
JKPqjmrHA9KcRf30oxI/ECoRsKzX1gDTSVmwRPcVEFbwdGEUEHW5J0DN1iskMNiGyq5IolyTxwfb
z12zU3Oilg/vsl9g0KgqUVVEd6N1z0NyPAusNquBnclXGv2lbHzSchHe2YToRMZhRUc9/af2QiNb
0ZC0svJkHaUKqTHOXeU6RTzMCLq4T84yDizFDsOYg+su30S+4GOXzLqmp+iDQ5baxBuyBHoiKhOH
Tes976C6Pk4qq7MMICzpxid1vE2ZvvShTrAnjOF90QWNAlc5d4V+r1Z6Vo9T++KLuiUPHG6+Nl0J
HJaObC52e59ip04NZvpb1hwuttKzZYdqVw049e2q+eRVYKVZY173113F63K+dsHyTRhB+rQpgrsU
HYMxDBdiRLvyQMvunYtr+0ns57EDe+ByTUMwnRX9XexCMO5xeRdK+xcxWmJFHXDoBcZS2CGJV5Uf
UK7Gtim8KBeRbg5H7qd38TVABDFuBvbFNmi4YlzIS0ltNxNbFsRry29W58WNdtHMiKlM+x9yNb1X
SLqf9ecuPRpOrQowxEpfUyvTfr31GWMknmaMoKslXLugEZOy3eecQw5DpuwLGhZPcEZOMnyacba5
0nCib2s2wlk7fIkMyfYPnfKF04BlQWFEDbDdSSAOedyg5gaWNYTYVSu+/1pRNy2/BJLGCEMgaM62
x7yKY4PIF9hLMEtojlh3hKR9yxBiAxekeim8vBXW3bmIGBTMbICsOmrK5iwc4jPepabsnGJyI2c3
J91OmUIjPupZSnrxt3v9enl2FWXxllX816eVKWRUELT3Mm3Yp3TwJmosKF26MhRG4CaYo5gnJjF9
53g2hfX/GDhtphFC9dXhyYazc5N4+JLmz0pjQOx9MaHQSaHdE5kLlduts/e6053b4g9sYwKqp9sR
Tu/LD/opZjGBSWmjo/cYo5i1rWFxtzkzA5KCDW2ty50h5F4nmUOzBqzhQ8hjS7WP1UWvax1EKY7/
ACBZEGGtViXCdxaavjFvh5oBai8ZbxKb8pyp+Ffx0zgvGKoj6/ACkNdchBZNosXFmAkQnOCoup01
HKT3u/1YFAy6AtjU7vnPn4xQ4JVlzFAAobIAqdSnSNeUMdFHZptaWPo1KdXcpO6EZgIphvw9HE71
aNHW2mu0h4BCPfDQjYom5c64xJSUL3p6ZxIkR7lwfZIr0vEObr2TOpPnptLXLZsaAUDDeoBwtSty
XVU0oNTJtH37hdoNCWPkAC/c2zb1GUssFhOGOooGfseYNxTy6ITKts2OGCvhXJO2M7k09d8OacVa
g7pkoygK4I6hbdBKcJzW/vuC2OiC8K9hOE493ekw4bjAs8fdgIw9GNwD6u1jzbCCVkXHEB4wV3s7
esfGNHuI0DMql2I3j4pcHfGUtn89yIAFSbn2lmIiAy47Z+rJF45HxiuwfQiid9Y5Fd02sOFr4t4T
i/whNONXZoQ5yP4SFvRNO4a4N65bSEyiumo0Ajn4DHpGSOUQiIfkR52xQIZ+oj4AgJ9dIFOT82cN
CwTfuTu51W3acnodFF5H3CmL0HmCQijZQQdqxb5mIXnwzDGm0bsVYGtkXoT4rXrrTudj/mv9wp7l
BiwHxyC17Ny3yHAwhWImQHRRv6Zv1VbwMZxzW3HqjZ+WHoBt7UIFNT5TEj2HYjbK0EZUltMTpWK6
TR3ZvHkRvi+7Iovb1wPB0v6efU6zNAB0yBibar41evRNP/Uoeeteb+T6/5oi1tw+3tJO42Eh3msg
6Zye1gb365U7j9WMls6AOQS7qDQc1dJPSdBckWd1YAAdd0Dvv6mrFSpL0RdFW1Nkotmc1AjjiRQz
s4IPWVP7VbE4Y4P2oObJ3ozD3hoPrhIL7/ba2a22425KJ4fCiKltRCEJLTfjycjh5Gp33w8LpS/t
WergH76Xe7qlcs+rrW3Qpcnfghdg5B21XJ8lEbfzxx0ll+23Ex432LlmkZ8DUN0HUeiRM8bu7Jlu
3uFucVnVGfcEv481W2YXccWgegmGkp6VP4Wfks1Hrt0wGwVSz1hIlWU1vkz/IuKaGi6ERq78APNL
I4QDSSgkHCA2Rf3WmbNlQ/8I1RC2PamWRh14y5eaazOEd3qabrkCwOpe2v+bcNg170B7oivfcG/y
Q27zwViNwCxEM8rWimC7ZarmJ2NT20Y2o0FE8TdvD4KjkFHdt9xRjKA7TG670uP19EzIjDhiujyi
/rjXR65YT4DS6IdR8U3yNMMlUWEpzeEw2LaoLrWgNolnWojx/Fh63o1w+/stiBm1kLiVD+kOK6ZR
cx2eu/kuU/dBrXaX/qTs/bFiD3rOFbmt0NG+h+G6z+x99eBo4ovQc3pZq2w9q8zwHS+JiORSORbt
fqzVNwkDYykIhusOH6SmCUp9UGwEXk/o4KKGXSPKs18A2GIgbrqxnge4b/q3RRhRLF1Du00N2zib
zAWpLRlZ1+PkcctIq3UUsZVR0N1MPTli5vYdWoM/3t1xq5xNiWDaLCij4DEbVo+KciiXwM6A1Q1G
wPLYMu/5ltQjFPSqeqHUG2GmIUsavTTLwq8TvjRKF1kmZDY9cP5Yi8MrAHYgK9cAkVlmg3DbOIT9
cdft+I0UtBgzTNPtXPdpTAWAUKjx5LuIDtFHALNlyVTXy+lhWDdtLKKp3GVGLb7zvc5/sVTDHnFh
1bTnKSYwRbXb4ejGh3OZX1lwawa8t160T+0ZrchZgv9Ppw34AEXO8Reh3mAXOszoTI6lr2LwP3C/
eiMc4sEGtIGQT5bwHKuM/U5njKMxUddxCXQe6DLQX/I2ZekU3ubqSksnLVStuyPmTTCfir9y/5Px
dC3n2OOxG0nSugwlEkrXbLInfRGNhzUnsMnIh9I4oD0pTF8wa2OD/yeNQMkoEymJtDt5SwwHVicC
TnQu8F2N8Gn9cyYl4vT/eOuPV6djU0dh+4UTLxY60XR/SHNE80Z7DTsJfVjyTHBxHB00qVc52oj1
C+vrVUf6Ki6I4MtwdZcxBfUPeRgKqaZzY+zpxcGj75zPs33Z7g5E3WPboWPOMTQqSNjAlE+iUKs9
ujevXnBaE6yse62BGzBuq4Zp9bRKr9ySkyXaV7D5dugAMKOH2FsikMXV+soBTreLqgXxPBmkgK1T
RWbkwZEQd6I+Qxnac/JxgYQJFeTHwiLT/OOXxkBvN1LPb3rOEx2fhFwPLkcSgebJzuuQ3dTsCAbY
3rMwSsid5FkhoYNKo/FYV4CDu4HSsFXaDFrNj2CNpuCDFu3A4rxPjRS//Alw1zK9zvcbv6XDMXNW
E3NM/qy7JtirJzSNiTiu8eVLkPHQkSDQsXerBALkY6MwKMBrHl5+1VihrRTCJ147C+tBM+r4wtIi
P/OPCEZnqRdtpse1gggJH9zsJpy8oqH8q5324HXBGDOGjgCLiP+3DdAITjX71lWkFv9KSc5ZMoLo
ZIUrm3gVSTHBFC5Ec7jMchwa6qrSsLQF94KxQQDM2swKYSR3W/Jlvju6V+2WnwpfrOf9K7FJcdnN
P+d8btHrYQ+VFRnuro1CBaPw1RGa7C7BwettJf8g5oHYg2WjMvGg8vlbsVr8ENcE7EEPFy8PFZWt
KPPobcdoVGa02zIDvlOY/PuUbDFn1smc6ey+fM+3KLU+tlaQA/ilMilPiYH4x5/sw9RI6r70UNx9
g7C/PEMqWj9TUSUilFWM2tvDfGwAjhtNWtjPDsP5w6BzJ5BGiwrQgxe0+0JHPb1H61C+fcOuP374
y2wdTuohEFxiSyFSMcMJJj9hw6ItFygSNlOvRzOt/H9kcle0C4Xxi0qsymgcwFLIG94000d44fvu
cLAnrLryK558Q2mg2LpAaSWBtQGfdZbRazQDrXOav0fr0PWi48fdwMAJQSUdjmrpeVqL4DdJBTLK
5w27hzMRwyICzFbVWLUw5nDGFnrt5W1nQlhMwEkItiFtdpLgxWXZ5fr3eeAfF2tRnRpIwmjFDFMT
4DZjB+wLimz0nV1WQ+nY92cFsk7En/b5v+NlS0A3X7Ho74cmKP7Cc4GsxIZWmAyKV4QbIQPTqA4s
SD5TogrENB6bWY80M0rzsolX/JY7WkFhFXPf27x1zLmnbaMHZxNMm9pibopSU8zRaMT3aVJNlq8k
FinFCrLU3KT4oFoehtQgTxlcZIBra1aqY2cjLwnXJsPE+ON9Y5gwCBZS+CJlPOUlV7UhXF2zjFBN
/CSA83ixDVX2pKpVuMFGF5cKkfh3r7/6lYRZlrbQSX6ZoKP4YAakWKO56DYAzWgO/UaXrCoX2XBf
+Ux3844cjI3kf2oqMgw5lMB55XD5iwKDVwAmbCQ29NXLEnVv2kerk6ZYW5fBLLtq5RM+mCqROkgH
mTy5g23y1ZCvYQr53ZeGSgNWx/5XT6JEc3IIl0Iat4qkQIrstDHGJiQj1a6usG4Xgc+uKUxY/66+
PnasXtK+DKM65Ko/EslpBDwB3Pv/xsOla/jjV6ty3TgJYeCLOa/ndUXUNWMjqrWJaxxiFpKPwbpI
U2hzj+8qr+g1mGgDH0zjkjJ0oYPTuEUBR8ThTmfuOFx4K+h0DNPmHfNHI9pK0UVppYFLuLPh0t6/
qE3oQ+WUJhzF/fbB2LKyn0j/4wfS2W+Z1Zf6wp8LQB3maQUiqNMj5wDT8w5xQZfoVO/5uw5Nj2tM
7dKT/ywS7bbqmMtYA51CI+9s8JT8DHRU/cdiD95Vh8RkZjyIXl3IIprsNdBVgh8ZYOGKcIMhJvzl
T5usc6SdXuGmH//eD49zOoZ5EQRkg3GwA0Lnhb/GxJdoy0VUGHqwbvskCd6+03C8+LkBhBe6NCqu
H0MepaBjAmfCOAQn+Ihgtu0cxERFll4dzuMg4GignGH0aQvQMIMW1NOwSP0BhwkNYpjcZzZeqI/1
QBaxpuEi2yOfdGO6HvScHi7CbhAsmQlxS45CzD07VPJEc1KwO/aDgSJ6POsme0R/17gVZwUdLvhl
3HwwLHm/nNrQOu2fh+Teydj7Q4I0ofHfkAh19j9GTchX0JqiLFQtDRZkMZJ1V/d7rw/1JpfacqR9
Xo3S+6XgwHAs2+pLWpCvYDKIEOcsXEWuC9Ps/AV/AtUsFyHI6300TeDHILqyI43vAXiYGxag77wq
U8/3upq3IpVFLg1s/zJ1S5lDjzZoJeJku9YFMOtHx5X7T+x8kF7T1g0RR55dsBasCUojYFXRjSu2
UyUlLPQQLa/d4GA/aDYwl2SqQHrm3vTw4p9iEtFVmtAN/V59hn6go9aamFJHKa/FEmy+UUlSM8tU
lFquSogqspOCnkNln1ST7EAN9+Jf+P4tNhkgEcfrS5n/lNb9frc9C28QpOA1oyqqgPM/x0YIubH4
6xNVKuBzu7swoDmjbowSbmR9UFdvLXwp/okCLpcREeACgV8wm8DHGWXEScBfV6it1nU/Gel3PsGk
7tO/yNIuX4rio2TFmbrdOGKR0MSO78ZhZV3oKxWC7pHZHMe/bU4NPkfvZqZpu9XLlMec7JQX/KP9
hXYOBN4Jk4Iph2JK9CMBapWzTfEbvLIunZ0Xuz+rOF1RyPGaecX075xspFavkGU/1Yr3S4EZkgZz
Xi4qxQX/OjbPQgZNZ8DfUNgohueHaZ0rOT6P0+IBNoe1Q4mX0WHI57vhj8fAfrD8jn/1R5/JjAD3
7DNdGatmc4qApOKFPoz85lW4Mpn3H50ivkWOOMWaR0LjL+Jbwye/hNeInZ9Pfyh2WoZoP3kFFdrz
gFkSmy4iwXuK5G+Jv3nynXD38QjjHTaeNpzkb85SlFusUiptwZDnXGN0q5zdAIdlx+aFDXJJI97U
B0tIw5YtsPa7uWPd6bJv7351XD/FkXPQcx6APYBtnxenAdPhxto5uoO0RYgGBGRS8PsOhsxmKSBU
JnTNAZtmUyiw29pZ+xHbTqFwvBt5g+JGBmIaqFB6sd98zRpdZQwaKXA1vvtKoA==
`pragma protect end_protected
