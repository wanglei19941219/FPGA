library verilog;
use verilog.vl_types.all;
entity ctrl_top_tb is
end ctrl_top_tb;
