// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:42:08 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sziNqyyQ7JkkUZ6hL2Q4fI0hxroZIG1uf69Qp3bScwo2fDpHBL3aQd632u9mD2JY
b772YHtHiFrLwEaQvIa2Xds0I0DHotZ0Qz2XmqMFLp4puAhqQfS/WOR8XWkykHKX
RinfM/cR3/GCscNO77nxqw8PI2MXq9MvRS9kyKzvpP0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6624)
ZUm/118ERrZiBIckngHCDKV03nyd2S7gesQp4pYG2xOkwG9KX835nBK1e9y5qaGX
fL9qXdU98L/OGdF0oWiWGgFQoKCoGPVJuvfWdaSVm+QIKhCRv8d1FHI8PHuPuKXS
cxPol/+fmd2dlrWLoX0BX+g/cxze6UD1m0hJqz1X4/CDaLbqTwR2H0DNOwAmFPQu
GoyQe7uaZlE/rkT42Gg1S4LZ9V/YeeYctDZ3xd1H94hBLGkq7vGkzzPl/nPGroSI
6pqZDKlEfG+UI0EL368P0Wl0gHZiiHpFfcThVWwaV0iam+6gxl2z22ml2SBUB/7I
VCVpxTgfyNHCKJFsWLZdCmofn/AiWFkPjfAEqKa/3v/cimZxcWOWlIl8M9YYBwfP
z1sp1WjYKl07X+auoJHRxtNwQhUmLY8fUXATy4JXMIRjj+5BXIY3mIbwkm91Y3w9
R3dMplinpMfrnPaUfwCJcyLdQLUvM5WT7RB4vGof86DwrCmb07dZhSKGit2qGeGu
d0esiaag/BJBct5B3xwBf035YNIxruldRNjdk2HXwq8xU/belVfySa82EM6ctscE
nXjXxcOU0oO7vUqJfTWQIK0YfUsXGasGEnfVc2kkEtyXO00dn3+hsDRSDjf2n0SK
bp6gdR756ifXTNZbUVVnlhaI3thJERWHpiaie/t5uf0BaSWx9C9AOOS5vfoCgCOi
aJR1M5t71SFtds/s8HQtDLKUGnaaEtYqCPuWdeWR19PX8FHeDhm433C4rHm68Ey5
5dxWi3AU7Ah/+ph55FIAcNNioXQJI4/p+oSqdbfe1D0FVs0FWk4jObhhvullo5bC
L4zfUxSdaUs4eSHWY868QyX8XHujLySbc1gCO7WZvWA94+KSb2QMlxW1cqv2FS3K
YpZOg8Jd3c/uSIeuSc9G+1I3upI/na0X3l/DfhIb87V7sflVRNguUdTbydjpDJ2r
mGwJBfleIwwRmOtQ3+oJY5PA6S/LM5FlrsMv9wGTLzxmIlWe6J+BmM3JSYCGNOlV
AchgGPekF8bwfWXF6i4XIH1WmMLb+Fr4+9q1O33Mt8Q1v64SAcoC1g3jWH+qivyN
MXZJSm7YIbiQVHeMfz0vU6L6Cx6FO5ORam0NLmWpIBKT54unDZJTct8skmRIMKwq
j4RjacjL+oVOPciCPSTl8vdR+0jIg3tJyyadfpU1BBOr0ACrUhjIfmi7SLO7eeSt
Fsxm2Xv959jlmgpqRhrxYTI22PUG01O+Uqz8T1TeDRnXFYxXyL9Lk7Fn7JXWCWWK
FpmoFxzN8jkzZPa/rPPSX0d1aMOf1+j+BzYfLNvHZsiR7hd9A7zDpWgVkYwg2+q1
ckVZj2tcPrYk+fjSpLsTDHblbh9cMtZbyj9sNvGKC7juIZUYlIjLzUeiYAKJFI5M
EH/0wIQxTF5xxSuibJis43G/WRkn1dUAdooZqcrozavKGN5nnEonsGY5P2gHqvX1
rngtfm6wsLO/DfW9ntBkxqbBIJjZyhMm0JZwALNXkQyXvnsk+oRzEHuN/PDjh97/
qesOmakO41yKefhqsL60h7J6q61JkSHG6W5kIbelxJ4Gbe64472TLnwaTUIbTOVc
qQ+aQWvZKmJ0Rom20x5EKW1b/gVHnF6q7jVPFzukfHc53VFZm1G9H3eBGDoM1NBS
V+KVREXmrOF4hNUfHyhil7aQ/P1u1jG6O/tBGiAeip7ULQLFCFS8u6/lm2kW5A4g
zqdlTsTQeL9TU/z33dVqdw5A1BN1O+p4whpviVb35MisGBBXnRQ+DocnniR3Iwes
Fq59NyKBRlWomTmZTommAGCo/RlqQxcpTsnm6l+YtXa0/vVtXibQHQ95xSXUGJm/
iR5vY9F3I8eRsGKfFUGYXtqgthibsE/uTJjuLsKZ2IDxUMD3sEM26NLBL8gCcFuu
mDI6fBL49oM2Sc4iQjpn1Mx5ryOHAGEf1HJI01czUZSc8P5V8gruDmqnQhCAzlaa
/DJVLSELb/zUXuB0jMqXnSccz5wY0+Otu2V8Qz4s2ylNKqONelMUEQB+IvKLfekS
8gAbgEH1idgnWRL+z1D4R60ZgCygk0ckMJydo+MVUCGpzBG8jNDpgWb4YvZMB0oO
F00AHyWHuDmptgRUfbBCHWbVihgPcSXzrP6ztMKKV0E/8zHA706p5dEa5LSb99TO
CQ1Zh9+3yI2hqFR1mhs5X+2rdE9VkvDNIN+DDMcx6DgvKoDGoSbplii4LZ7C/kgw
xxWTidxGASQCGzkwlrxy85O42NQ13oq6ihFmUyyWsCgRmbTZfQre6JkzSgEcc+hr
0TUZbDAkY8T+FNpZT+hcmzuSayYSOZRKKJGwjt6spfCy/M8iG3pFQ227PCxnT6OV
RcZyEs1clPE/K1tDuRavMA6tEruWoLWd0f2lh/392iRC4oytwE6VpUtCt4jjdQ/8
DxeVQNDibAacmoLQuAEjs8Rz9b2n0xklqysGBkt32DaIVivuGG9YXA9J2PPfEjXJ
h6bKS3DM3uF5DbKQlsMY5Qmhh7jW7O/XKAgQ34QFIRgCfBazTWftDVznVrd9cJbO
+Zpe2FuqwXX3mSoy70cBy+pJxgdH9wu/Eaw9NuFB7xDiYb1AVDhbMGlkgv1Z9uIa
itxhKP/XANSrU8B4FuhoHngvDiWCRYL1v4CyvQ9RyVONDtMNvbtpJcpItaEvMDM+
n2J1dNmg6N0DEHbMb55avKKz1mNWplF1lL+LuTnFsFNk5dzHIK602DBNUEwEW44B
Uf/UkzGUJYI2R70ikdwvxe93VGgoRzB1s6mKthxtXaVcqE/L9tWYYclet7TO5oYc
EevJky25IodC7kg4vtFmIg73YzgYwr2LnBLf1nhK9yw9ERQkbAkaq9G5COaTR4nC
FXt2S+SZiHUCmcbQwFx0BhkM/YJ8EhKEzHcaybn6L00eNVYy+FHQUqWKbj2DMzpJ
gYieqLswZJcyYmvicJhAFBUfDKWqxeozbg1s4fI9M2oqZEdVB7wbnCHWCaK6gLnr
XrbHwwGAfXJ3yR0AZg5D6xM3B22OPpDAdqkhqq9kFoRTWTp/1OZ/J9rCJUMNyPcE
BHYHw9hVeGPC7sOgAGHatIXD1xtaPgDAjoeVjjley9hbTMIjKAS3PuZxm7BIb45U
F9XFsVfTNZs8pZkMCYAEdAOT263yQlBIrqYLDON9Apg+8dIMf7hL28GdtW1ObbqI
QlAPmP2xRVORaHBOMal3sJoJMnNE3mDdxnwo7zcG0yyT+D2ggfyMcQVI2GpIZYN5
Zy3JaB2+niO313Y28rCffXvMR9BW4CP+sFopJIGnJXh0JVC0E+jCh/OWMLbQ4mrf
KoUpTCv+izDsUHEgPAZlIcqEacp25sFOQIuvcxDHo2s9J6vyzerefGUBw3eLTNM2
UXNw09fpikb3LwZNFvV5AEqi9RrVyQAyBuV1G1sE1HtZ/6PM+fPWvy4DsAhIkjWe
HNhvoVPq6MHDLwV0Xe82F768XBcFtqjN7OGCo9jmgwJS5Q7YXZkpibcYHf4frJ72
/I8Ekl12pfRhgKlrtWGefa1vvd2PLgYJZw6Nlk+5IRrwc/VhqEdRlP6EiziJAvsa
Z+WXiG82zqgnBqvceEDjp/7mcBKnQI52g1pfUQ/6Ok90h74qQfAR45AG600eGde+
oa6IrGdW2BTF9PHOAtIpU88a9Y2JcUhxzXGtU+Opt8gAK5TW01Fp3por0jaEijS7
5lriTknsXE+JvbDLuiVnPE+zSiA0SUf8n4Ke23OLpJn6OVyLUqvV0V6CNnT9gcxV
xT36S8S0c1cNcN4dX3d2/emLq8LlJpwbYaqAioe4A/x07x0F+BcPhbs0hBXIzOXj
GfzFtSXuBXHj+RCgTknK6gBRFzAFnzUBCU+nrl/QTqWBRzxKX4hGw4D4/LN8apM9
75tv0Xt521obvlwCfY5NeoFKc8AButw4Abfp612k6vS6sOVhElmMwQm68BSZWk0W
sIoK28AeFXMtTwCryRDvs2eaPL23lXpCMoPtWaKuim0O/xzrnM8KYpRogIMjazs5
QluaDwGUf9j92ufnIoh+8x1ueHurBV1deaqNhyslGKWzeMOXumowzvMpAyW/NRH9
irnKJn+ps8dWHdCTR1KfMR5/LB8maoOfl+Bc6R5aj8sL9/zvMkNtU6CmY3bBzyKJ
jjpgiApxXV+9XBghsfATLRKT96mA0Mg8LOhmmnQG3ZN/e6RQLHBmpRo932ghZwdn
8fjC+JPrHiEUIPdv2x3Jusfcry1khiVdAgLHritMi2TzbEUo710LwfOoqWKywJRY
pLOSo2SE4FQ1TwbFOWkL6YjWkLNrCMphPf3ggc/FLQcBSMkQS3rItprMvkm4yg3Q
4t+jJ9lqoXDR1QkRDDPbs45JzOfZyPfyzVsObzpy/jjfCk2pnsf6X93ig7j489yK
q/Fv0H9LeqtxYJtSd4zzKEMo4qHs8XL9orB362Em3+snReIT7YUkvCLkSFb4pnto
qtjDq9OFWiHqymwaFu/b93LvsxcMt5cjxYGYBYDC0siiUMI2BLna3S12AZMAjq/R
mEepdbRxn4gpcLc2N4C1U3BXL2r9beckutWwfWzP0j4xtqlrwYKLyBOrAvuskNsY
oAKbPLcAUMnnOzzrYDWuAKZI2lJ2dreARcf4esCexQUDrcBmLbPcpWzANcTUWWDf
JKRjaSZ/fAgALKQ19WLOp0JfwwmDnAIRjrZeGH9NTQjC8g0F7PrpbKoQ49Eq0nmm
r6xfHRJC41urIZ0M4C6enxMMouy2UmKdNlXmYMMVykaIeYGSbXQlN9STRBDSmz8m
jJl/zzmePGI7pDWUKcQ9vqFpFIlZflOJfQCagApNsoqh28Xee7yMjA/PcD0NA9cR
FeqMfS54+C7bAvPuxBiD0ux/Y54vybxfU+rvEh2RteNvPTLi1TplTWtMNZooFSpb
dShf7KTrEPlfwbs91+gYQueJQjZq4Dheuw3TBisBlFDg85QZ98FUQEqMSgQUt7kI
vSGy0ckQOWGXOFxRCCnCHN+fOkbbeEC3gg6yzFr9TN3vlj/V1EBaPwFhi6NJYp8a
9yTPHJBFFJPyCiGPu7TrzSTciVL3+W13C8Z2c5HXDCxxpc6neb3ykY86xKQhbmRR
MlmjKoo7rPfhDqjRXX2j8coPmiqXeREspa0qSXLADOstw0wnz6WtwqA88S3hTNBp
wqn0sXBKkoh2VH2OlFZ2Tp3cPe33MtZZLCeKtVdw/a4FdiKwopUy5jIqtizt/sjE
NhG0PcUDzATlg2LwWN8Wa+IBpgznBZDd9NuE45z8hU/AEPsvCqIQLKplEZLafnVy
IHfSinOAESNVwi6KLdGAsstWeLNJ8y1xjjPM/0RpUNVmXM30DSKCax4I0NohMI9+
GO1HcnCTb72eqMtCzkEjJj+c/vhO5/PQXgTM+xSPd4JCKEpBjGUgwWUkfF00wgVu
ecpd13n1dpOmWxvF7ADySnl6oH4na0hzn+6LG4D1/UX8RANgVLt+WqPjKz0MaJ/U
T7ekffOEovCUD7uGZqNX1U4cQaIXnVylxgBC2zZFitV56ikvaVYCzGenY/GBPHRQ
R2JDyfhu165IGP7m419EtOP+zX7nj9ziGcGlGOTyG95WOYCzMN/2Kj4aGGrjRVio
lhw0w++DYyyWqbj36JTXWaO1KJ3gB1X7t7uC1tTnsIJN9lnKVR/zrx/1JHUC7L0R
tgiDtq8MgJPcI32igk22TWwHBePpHRxFPu+lVM8oF+scWNdw6+3IO71tqY85lTS5
A14PYOobh+Fs2f8FX7Hb11zYNkAwjI2KsDdcCu+pCZB8b9qBPVDDJRwJ1P1vQhLW
IrP2BWtxssAnJ8ogT1J9VsfcrbS7471jdvOEH/WoTfp3GQhq6dThhGwbbkxIjeat
MqF055VFuflhjD7V8behInkiHLk9RHiGr89QB1BnO7Vn1NntJWUe/InMxuypjQVq
k9MCKKW1ypbJEPfw8xfrFUkRiPHIQLWCWQNAD9Ywiv2zOE8LC0+bSp/ErIQ4H6bK
lBKbUeGasENNTpRunEGON682JsZTu/Po4upFpVjUH8pAUcFHIWOonQkk6QYdErar
KAT8mGf9qwgeEWhVmppnbfEjAsIhPuffNiZAy8upLcZyhJvg9ICbrQwoSjAMu4TN
uXbxJsQe81E1tyqsjpPOWfKxn3o9ATOOBcgtWyCTg9hrvdIPcCbR6OonvMh/wlbR
n7YUC54c3UXhih0bD/jfqBfuntEbhH6RkQwhlUn9TnzBzOkfCfIccjuqX92BRKJf
1hhJQSoOzr1noO2PgDxHS+S1xL+NkQAtwxnxnLbC/67CYj0pHVQs1uRNZEwhjtzD
VToFegCQXSDOfi3o6/EoYg3wkgVFXzi9KzDtk0fbzGY9xdjtG5Ai1NM9MT49ESMX
xRIwGhLo77XAgJI4eNfeDml5T7xtDObztpY4skEJMB/ZAlJRkZdT5iZyszY1ND1Q
SEfxXIb9LkplfUi00chwc5rDfEQQxhCSlHZx1eb/0ibhISNB2YoIjRs0VaFVQ9J8
L6GmqTVHtz0Bqa4v+GEx4TYcg2rD4MkSACCu+BcZPxN7bPogja4izIJzmyc7C+SB
ox0+JLaU2mB4gpow+pA3I7NDIqqRq97JhnO4ma+SiagcY2zUYzuaYywoLVsahMYL
W+2zh1m/4Dfr+WPQdFe4iRqRo9mI6Sl6e/rMRpZILFr36tLQEtxiDB8m6pdkmGLj
hXhKtyVDq9ScTuuPfHNBs0buTlx9s0NCYkrGyDGRDb2qyRJDwMH1Ys9456l0Evu6
6vTJ4JnQZrfp7uEK8rmRaOHCnUMTknVawbKBMyTUpA3qVL8jC77SST0LabwRkTMk
vQ4VleGTsvwkl0IQkRxpcrj9anlh/r9rcB28V/omY3x0uEg4lMnnEnVadDRm62fE
i9gKsHSFiWdvTiY1MCu/8mmjUam7sx9HXBIFKEQ3lxWpja9w/nyYFUFIlUEbzJRz
+qnY3My7Ad3UcKM6EM0Q+dMGbLwBA9hKf9rzO2PTP0gQK0dhVKr6NQukQmEUx5ly
Z+/0YgVN3MSQdzm0uL7bk0N8JQd0tRskNI+faPKkcAhraxls8pHCz1KFQvoU7nyz
Mt1pXnEbJoSgmB9D9tAR65G+ShYm+o6LpClL++wEGTua9011ruk6hL38PR2r8QSh
ohll3sYJ3EVm5RtIXSFABxglYiplXH/BQ1h9ZOFzl1Bo6blFmbJxf2dlRbn5JBxs
l2KG3SGi12JFxI7HlyKR4fh46qOaKInqXzCSzA8R3jaMxJSsV1vFcLStkL2s5v56
8/+sVMeiZreghJe9dgG4enEpX7Xs/nBDWJrwYvYTt0ICcHavYAiUqisWNurnxrlm
nFbHd+u/MrDgIefidlUVmd1n6svdbhmsdqsB+PU+IPkJnN4BVH7MO6HGNK2V2ZH5
DIe8fB+gYpHyTwBgZBLdmL7MCdf83mxew5ySseRZYsTPwFfcYu8bjAG7ECiURHAl
pnrn0kIlEQKFQYc1OiDgeCI9IUpCFeAz4+BVte/nyWVQwHRBtDCVeNuUViDH634m
oavNQIoLBuE/KAh6u5kjzxyLEMR3hbTcCbF1ybjqeL/t8Wlqz3wm1Wr0otopeg98
LcjnRNf3DMLKHTR6fYFzvskVE3wF3BMZ95RFiyjpio6E502xSq80enB74B8RZpIc
peRVcfqwE7u5M0jMKUjKD7DIv3Gheuo4syYT9GJpkax3Yx6otXDdtKrL/Xe1WzWs
tP+IhlqAS+zkm+/ipUTHuTwqM17FsG1WJ8yAtPHjtYbBaacqaibJqU72D1Cf67SC
92ZyKs6uLyIjzcIqVm9oY4KVBip/1pkYJ7MKUsRcXXR1kEXuc8REukvZ/IkGGxE5
gQD7kNekJFTtCjrhnHN4rGlqiW2+sPdiAvzZNjoq9z3havSBSsjvIv1sdUwuGlFL
0NHQlrOQ9fUqfXGTaGpoJJvOfSPeI17Pa7m/6y6whZmsNQH7qJw8+4PPOF2+QWQe
AhJTeqA+r9kWaXz6AFb5Zq9ye9TAYNsvrVGCMDrJxgWbo68K0BHHOryhyVnivVIN
/j5/KCBb2RXXVQyfEhaFgAHrp17Ea1KUVPDWLVZ+ZpVadChO5hm2HMierC5TBx35
kiwqrVF3d+aBTDyWqdQOAVy9qiNAmyWaN/2uubzF/U3+NpDg2cENuCOZGzLjQ/2N
rSRyHYhKcsv35Cu5Z0A2OLVKRI5TyNr4pQM34MUuVnmCXwI3YdHg8H+M1n1ckXp2
tm6j9GOLyoO11kNcn8EoglyuWWo1oVs90xDj7j6c9RXzT/6eagB8/MRc27TQuIH+
+Q8nSB/X3LEEgmQyyFsU+nZnCTHgBFCe/OBKtvmd+n/40xKzC7wLQqJ6ZwVBstc0
oE0abYgyQUONrW+farOjUaIx1SRsbg9b+mMxPkPWEN1zPug2QRdJbyNLc9UhG/I2
Ne7ReJpH9x1sT6lFkgDkGcLlQvh9I19j36WMuYeuDUxDEdICdv5sjabLrryUQ8IU
FrbXaK3flqm0q/uCABO3ARo68Ru43HiIoaU2DGWNuKhzDgms3OURYnYuw0hZ27zC
rH96EyvGj2mCz4uXdUgDkh6DKL7tq1pfEx6okuyf+oR3XpX8Cv+1kDGieic3tlut
KoNH3awO3KnRydkhWcgoCOsAXirQMOe71dOzPhllFhqH2cRRW7fp64tQEHcxUI4H
lyJQ2tuL5v/mdK8aF/j1gwqhSeCu4r5W4wA4nxPt7CgB4C1mU2WuZRb730AViQ9y
qZZtYW6Lo85b8MrRFwqS96iRZa99RrQAUHYg010RpKKB5NHHQJ+rhNcHAblUPPzX
`pragma protect end_protected
