// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
EKZUFAmcaPTq25DD55UL8QmlPKpVlH65R/9MR92ToZSTcs7X3znHXJW6K0Ij1i/DQkNt8lmmp4RC
paVHZJVvMEsEFNnYqI+aBlX81/Jmwr5r4YPFGK6SRnIcVGTLs+Ux/RuCWueF8zD/WRAiO+GY3OU5
n8YW8PZWiG5//SQ5PKzD0zHhI/9rflGR4nbcaFfbEggQncizJC5PELlPHv/gj0BfIC3Ax+tQH6Jc
jjlvaAXBvOO3bRFuRcl9C69zAVPnUFOAS1kqCeQqa+FZ7pkYRF1uWUWmvcmjD021itM/+9LTYU12
sqXy1LmuK/JRnhYMulXu6lxukNRIBMeCd+9ZmA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Yke0yJgRQ4WrFjwgCu19ZYyxRGSdPTBcxUp4H22ZlNmzT/G7FBaL28ySVCyqYPojLOa8hpvc1ah3
UwJQlio1A0TdQ93ooOvfOtIiWREDr2isqqP9DBJX3bnX5oU6WwKZ8NPJaxzgs0URuBUmZGSxKGir
mszO+fB23lt78wRDrZVJTdT7SoJ2e4LUf/p6p6PQZGyxHBhRjGrPlz1G2wVxRIdPqxyVGyxckIfe
F/NpF2LJ/U6C4w9y8IJGdWxOex0DjalNePV7gCYS6XESKEQePna7cuy4xngwgTs2PU2JB91rCRuP
7kWB7FQSfGFi0mOYEotRSI+uNiLzGvv3Gv4r2jqHJ1o8oVatUYTZ2Pdh0QGTpV8vfG39y/MCjO7o
1lFnRO3nJA+jFt3YhUKqIzHNUvlqlHeCxfXgKnZpD2mo7xmaRcrBdAEekwUj6O3KVNghDcldH4Ry
836wAQBInllGL0zsDuu+BCjwvBjt4Sm66or/+hLqLmAfxEguOV7qlJVTvoOVloCVLUzHJ+5nOqpQ
sRs5YQnVkFZQIkdfcBG0sZ5DFI6nU5jWTLfwjxOC0vqoOyQMnDrPdJy8Ajx+Z9q3mXMS6jEySMcU
L6XeYn5vt3NKcw397KNJCQbFiGA7Ohtn3FmNhcXt6n/Urvia0PcRrS+R7jJeGFQIqvblPBfspRoU
3lLNEMDMCKh7KmMwZfW4yv8Io1byVMi+YVFcGk1/mOTSLnseup3SQIUpotJAES7MAUHI+4mTjMlU
5V4xHGbzJUwKMzRFv70TjrVIJPabNG4itzAqcbkec718IdiHQE9b2Okvfq2Zz5jAxm4SOmck4Cdu
ew+n7KjII6Z2BjTJ5Q0OBfws/F8OH2SJAAMzx6CRBgRKlxSR9Y8/tL/FkNr6s/VUr+1CqutGVQYh
mmxguujmy3VgzghCGUPiZQxYyLMHL6LnXzBbPT5OJ3Rteb8mg0GshhyGDwThxobhfKc24d5+k1cW
KDd3NwgRZ/jo+HU94Tashf3v21TgVM+WpkSUZrhrDK4HseVMoJMcT3jFpkCgG/nVlet43grbx8Qb
EY16k0hHkLDFp1aUhKvKGm5dY9R1frB7ceGGwYJRlsc3uAlS+XhNVb7S20rVOK0PWiX3O89xGAEA
+IKo9IswrEEd/B+HPUQxFVnz2ALd8uVm+0tzim6c/2ULDrX42JFnTX9Do33Jcnev8iX0Rnp9l8IH
UMz2zADr0CVfvBDBKsAC8MbCSn3yVv1aJIomFjNN4A2/dX+kgR3ZfAjIAft43vMybRKc6iZxbuRs
gRKasCdI2DaplrtuX8J5c+H6zKLksaV7lMP0zNbS3PLADO6TUCXV/SPi3Ux4uxVLK/SVyaGxpZai
18uHpZwM3EUz6XZZbU5wpVcgG7rDpmFBNT2AUbGSwAoAhzoKmtpImsGYKBTmmiHFz5cjqk3cMB3e
ak03mUF/NVLJHtzpM9lpGTfi0NiyfqsIgvCiC1GLOC2Z+h2HgNgAger9212mDQA4MzFOpgUgnEbS
nhaaV9bvdlDyHjkXPmOA0mUMr6f25iJf1EcqemgSrDlB+2w7FZe65cJiZ+cMuS4LZKd7J8LfE9KU
0WuuUXY4xdUYduaJDvwXlwXL0Ubn7JwaR79FoKhL//RgoYb352hM11MoL2F1M+e+EiDjBwLFjGql
GiR4pbAu8/37YmNrZvIIHzWDRJH1K/CuMGhTeg4ycacYe9D2V35C8b+KFPy5NkQ4mZoOq6t/qZU0
kK6tHe036laBcN29ayID8yr/gqTJ7iCC4kinezCkATyqzDOQALiQe8lwvJtd6Cm+g4erVf7VxVt6
nEgOYKZKwxm0FoCPX/2q8LwSn3FfW9amqmVb9poTldL6iBvfUanrZP624XEFrIethBF49qAsgxQP
1OJYH5bHbSoKMRBpeFZBVhKKbWMLbfsna/W74S3Dx8emMkICIS49gIvDt8uBdHH8czg3w6+NZ3ua
Hh55np143EmtHNv1i12v23xqwcJsYPEKKgE1xihLrV/lQzE1WUhblOXjiJS4n1B3uloBxCbJLzNU
HOzFykOqUrwZcPkdW+Rr+ga8sCT/yFOI4Z3pCtyqt6vVHepU1ZSxHtnl+I+Qz1rzcZ3dK4WrkRWv
F9Wm2hduFBRvQWBvvAyl38oKq8WFvlxTJxp6eoJwDUaoHQNHgDf/jC8s+BIDbXM7X+QafMup9Rno
xlvLCouICMVOWvAvW+SLlPdOTBXqr240zB0/8pJMkJ71xlRM/D98/YOyqJia7A7cbbp9idBRWRRu
u0neuhHPYOJ9BS7HREp3bnqbEcldQrR677M6EbR6mmKtCbKVZk0SHURaZz1blxIkqMRgcopwjUe4
8TfVqcIh4JKUmpRg/dda0nn1YDX5SNMMfj849ZzEvRRxW5BBsDfPZcUcsbwQbapCmDQXCou1vxKM
mCOxMx5RoSu1iDzd/RX6qCyRpVoa9oH1xH2Q+VIIT0GDKwgDuVOJCqMXZ/wbpDMkBjijKsvzF2Hs
JGDPKZt/meNNMk1uJx85bHCNwxJ+WJEsFp7Jqo/qRYTeuz305F16RnqHLPmNQR7sInywZfMc0iMs
TV1KkTRJoP8IaT+cCNx8Kz/6DOw0MGmcN3v9V8xyIX9XQEcKGyfE9eUfwYl+HlVTvn+0g+WqzhBJ
wm5vJCn3Yb6P8q/SzgU4uKiZTVkX1UyLCBaBNyzj9BD0Bi9N66xw8rtcYrDv2zjhtmsIMqqkm6YF
rm9kyZSNiChzWpFrcW/281g6F+EnRcMtU/d23B4TRqjudGz+s6l1XHk2gA2lP2S6H/b/0JP63ABb
aFEHSr2iHe8EwpJzUkyTWs0MptSbiMOTHEjbbkAv4vxKsvWGTaUwWQDkd3gHh11GeeIDSwbpWD40
24hZx77wg76lv+/AuwTu/shvJaKZWkDM4enS9qMQ3iKtNLlejN6r/1lXsjLgQ/gNZB/4VnMWy2PM
wUNMBb7nr04z9azE7GtI+zM2uI5HpVQyctqDOz0PU1PMPujpYF5mbyK9i0th3JJ8GQtU0oY5MXog
l/Qtuw6lrXNoXfHGn1A0wVjxbSZdvDK7xzvm0cTvSyN5fX66/51lM5YTFd0YDvxwJZ4JCv6P88c/
tE5BFZXUpsB5PoLH6CaW+uf2CDQ7XLn6UCbUSnkxQoE4tSFv3d/R+gZ+oaS1nrzx6a5TQfIBrqNa
RDABAp87/O2ecYjSXHt1G6Rk5xfxzMcBjzEGkJAZjcbhGofJSfoqUUb5Y9tXtTL+MzRUG+kPPVcq
dAjGec0DpdWtO4o8PLZvaQqB8NLNK0yfg5dd3kJCUyO0mgddDdusiMSDAKQcC/ehyry7uEHILA8a
zfMcCcjo7NrBkKhAMS9HEaVn69WP+6sRYRYHmkUNvJBgjRbTkkV1xYJVvPAeLimaArOTqigsrcyE
kIkR4r8CSTrRaFUdm/ZoJ3tneGDZOPSwIOqIlQLQpHquu/PQVM59+5K/5ljgD/DClGOPoaZvVxmf
bFc4rw93ck825XcarZUFsQZMeoqO6/xk2gV/xRgsSirgWfNKyHKuwDRTt2F/xwdOlwx5yQZuyLFO
qAkgcVv3nU/nvrdRqzRxhU0/CI5yim24p5MunJ4z40oyyx6X3sc0pV/+1Xbe2G+76qY9MXWPNqVb
Atm2RBc137crZjS9BjUxS+XNKhHZaEbciIMw0qWVXm3k/jjYtB3bhiQrk/cDEqQ4dWMbpBpdXFpZ
GUzWvxgHewgET9b72HarTMC1nH2Gw2edsN+8keHp0p+n2jRCfNiMndbxCPyxYTnAMHezjLqqs+vK
w5MetQiZjyoq80V/L1F7CU5BzpYVGtXm5dStgmkUCiWD3BKm7C5MEGc2Rt+uX1WnjmqI7II7ZH8x
mEf1FvDBdMnCtpNkRbmmgbv2oMwvylrX8IWvIMJ8gyhhql3kxj/F9aUe9fasC62CE7Rqwv8h3/ov
F5i5ZP0LWQE/QXMVmkdqRBR5wv5bE8DNKxk2FFkK/0oLNaUTeayNU8wp0J0TiX9WVuoItqW4BHGN
U6Q6NsLI3qvc5Gir0xmj+bXMvt2Umgm632VQochZEzdlOwwuuueFOA56t6gkqnhQYLzSgjcymKLo
nvaNrdIVaMQlyjsF+/7LFAPzy4I2CykkD24vjCkGbKrzGED/bEJYf3qgMovdxdWI6o7YhApgf6jV
7YiGZ1Ie+08341PNa/doFDankjNFqJsWR6m96ol6iVzH870W0cEYKIwpQhqxLdMPB/wbOBRKA4+u
I5HkIKZT+9hiSyShT5K/+hDrve9iqtlX5GykFKVrSf4igBbQGnHt8fdrTV5mlqYvdzllNOw6Tph8
VXexNBEau2kVwMVAbrHliU24ysj2AO9EtZ643wSzyiFrf/AOcDxk5cR8o48E8DZsGmWdGfoEkYkZ
3y3280VlZgQs5v7vu16PuQ6uhHr7gnLpUM13XO14leHvguC3AXF7AxMrMb471w1Si/gi1lOIvY/w
oJba/Rstl/FcAjZAQKA5AUNlai8BKLu7PyvJ2qVe9nIK13qAQbrGfkWfxhXA0LvDbGl0x+Vpac1T
FZWjOmDNXww8aOBx1qPeTAWe9sd9tsYE+Z9dQ0jxnPydXiuFZHFzlugkNVeirGPwjjQhLJuwyN5F
a7j2dWqyQ4blI0Sy/aMvu3k79cgYuMi2VXUnYfmzw0uZVZdkVoABp8EExQV5NItq3aru71XdSxhA
2BNLZduvP/orH+XjuOXBY1oJwk3H+oYxqp9jg/BTGs2CG4zYcLH9mI9FrdEDwvI6KRS5pcysSx36
bZpgHmUdNwa6SGwJtn9iGw/siQaRpuqW9ZoiIG76S52hKyiOqWFvKLB6KaPjgqEbQVhAJPSreK8n
fdlOctDJK9D8hkK7Hu74XH893lN862z/Q4g3ziePBn+QsR19xb1B8wJe2+L0s1anSh0j9yTq+/o7
0mO7ThqlUdhYdJmy3xRQljfgZq0v2vZSOogg/fvQ7NqkPblzvBQg36EdAWTr4MGXYqFD0g0s9ccF
3okvZtII9k745RMuJl0HGDYOJTxLyw8TWKSaCJXKxdCmSaLGVJmMHRCCHcAk9BiA2R+zu6wd7Je7
bRQqg1Fbxr93naGTuX6Wi0PQbepXXgydL7su9EWyUtvXHiVqtoP+safJqERYQYqcuegKegyr0wML
MGmCmd2TML+4rGaZmz2oJh+ufcBMm881+dJctTeEl1O7CWT5WttggjddBzrCF8VBKHKB3/oArB7F
eiuq2B/eedF3jRnpiXPiJFNFwFCL+Zpz119B9hxkp8b714gUKIN+BIt2OR7h3MLNhehh5VuUApi9
/NoN/arxuBU1m5+Bi6eDfKTMqLBwIAjVlXP+Yv+FmPTc1Izk3rN4H82dfILdybvUfRfsWY2Zg5Ce
AJJK2QXrygaaNvJuuC8eELJ40otdBaDJA+vTiHgkV9vT9Ymw6WUaHQOmfH5dwTprU5l6am/THEIz
vUVHAUNYkTFz7m17Gfhk1+ABSsKEgCHqjXlq92fzPEykytbBXa5fGpMuqO6ObQC99+uYvhAFy7ZA
01rFAVifEB8NjMMqWFge4oyxqXy9yjUujTk9NZ6UZhyWgPdNb/BRXQhYWR2QKlgONR+Fy7UDgfwE
wdsU7JF/rQ3jHOsJXROOk/rxET2ImfHBK3I4Q5VTKg0V/3+y2CaippBMwFonKC1JzGoltJFjpTzR
HpMwkTVy7YgCaaR45mdQ954LpQhSwzxBYBEFJ+UdRT0Mc1wrvz6n1zkG4PGQz7vOPKb/qQDmXWAY
7BB5UXMkj3ANHZKxzm+0Mx02dMh9qOJtJ3kwgt1wfDEIcrt1L6QaEqJM7jRVZdQboQEt7UUxDqi9
MWZLCLTKUEoRBrwUCbaeBMvrFYzrwI+EdeWt2H+e6FZAQJFYhj2emGucb9+F57bddf/aqMjQ0Gki
KOoyZSpdOvpOcczanlie96v/P9SYh79myoFy7fwOcTkpOLiXuUjtjLkCBFkGmT67m4GuQyGuEnb2
/sZgtHTLO10fnory/VxtfKfXovCha0lReMaDu1CVhwFi59oyVeHCh+KwrqnSFtCJ9/07gwG+UVq8
z9tBX+I54qxaGK8vCCR6xq7e7p6Yzj7PIoWNxp5W0BXIvakrFosxMQBSNOOUrOnE/oRpu/1+FZZ7
cYjzAZxBx5qdHnkqE0pegidSwrL13D2JaamQevJQPNPA/9tq3UwBhK0BdaD4W+ta4/D4kpd9KPLU
NI1ehQnh3TnuW1lJfBFDUxlzYHDizZyJepo0DB+85qpBPOdYFs0uQyv0olpEQywu96ATveDQjsm+
roRoX0tNSKjin9I2/BrhL6/yXd3ws304kucnKwxaEDtjm94ow3g30kyTlKHgLJPJstXTfvuRDpoP
PFIeUHxXH68eyDpU5CwzwyuUatAbIS3t2QhNWNpqRCCD5o+P/hkoGlUAUS+MZmIH1mczcouXAwsF
ej9pqpOW2Ipah5ZW+nqUR9SL+jU45zWNzdBwmHB1d+6Sh1q7mvkhyCY8jLfV3D4ZiL8iSJcw1Y1i
p9ypCP4WvANY3JoLeKAyEJDKZuvlpT6aHfq8fbe9nwayYYASaAp7xKBkTpeHK/C94o/jp8LaTCk/
lZCSp+vyfqsu6phgXPB7SqwKH8CJZpzlaKM8N5gNExVMJnya291MMqeZPDPmgmBQ0Spe2H2Ix4wD
/wTALqCxKe8Nxs5j4glI/C/vZe85e+tpTTaTeMq+62BUZnUyadYtWpaLCngD9ICXQK/WfeJm/RgT
tyvpWTb5NuujWnBHL/IuWc9sCbCKYfWYeNYqaRIr8sj/4f3RhuZI7CDaoSma2FL4DtclEEuL9hMA
Ft8DEZuPVp9D1EhKKWm11L/ymE/lRt9nHLImgvIjbbO6/c4Gpqz2vGMNk0JhjJV17ezI0NVW86H8
S2PlxACiPlyjDof5+uw8uLe7cdNKjlRakcpCDiXUNaRCziT1FrNZf8vt1eOmY0amyBNmFKjzKLml
wkIL/Cl2VJLOocSlvOCiWvqvRiw=
`pragma protect end_protected
