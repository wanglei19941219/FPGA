// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.0
// ALTERA_TIMESTAMP:Thu Apr 23 10:42:09 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gTLYqkHhipAVInRyvaLUplD20aw+hk+DI0zkcOxvCw2sZJFzIoqhZUF4ZwFmsSks
/uqwcy2KEiw3Jh5XQccNha55Is/lK/J8X/gSZtwFo1J9KB09p3AtvO8kyYLgFZuW
fFVt58OfGC7cUi2ZpShlvO/gPuV7oCH+pExqT0XGWmI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5360)
+vrFZgP/WU0YvAcM0eQnlWTywhvtGkJ+KvpjGAy9YFyKgOYrRm3UNqH6YooZNhDC
sO+K1jTfnyXoB3DzgBAucs76e0ocTt7vOf1UB4aWaJqRFbjs1BdRWHI3tlgSYOpK
M1VeKjfKt36XFvKgrLATOsRqiAbtYlxBpOYt1DnTwR4lz61FvNyraSiYm8mTeEwz
yhlxjB6Hdwivt7aKYxd8ThKu+mK/zIc9XkN1oXX+Zcak993KzfYNOQKGlXvmzLq6
AsobEXlHhj8vAp7WwJaBTabHjJ26n23XRYDm0VrNgVycTQtNHdqwyDFxIXmCb70t
i1f4z+nL3yNPr1/0MgXuImZigPJK2ypz4+DrYxP8jcatDhzTkcYu3cNUrfTvntRI
Pu13LEf5Il/RS9qpo1CEQJYdtQnUMsrXWkDeak2hr57pkHGcBzVpt4g0OSyIOa9N
TBp6lE7+hmIrIuLw/rYrIhgq1u60CofkYe92aV1lUbmFE0nLV3hf+Gk/wwFKZHoA
5z9FW5sgxkAqUXGVntb5jPgJjYllnYeKFso5j9WjCRq0ecvjIC5wSq5ySkT8pf/T
PFZtk3Yr/i7Lq/yXNqH0xAKFqH2Z96z3M3rcid5nlxc+O/srIPkwhrRGksRubrzN
LDONJHD0Mwz+Jx4n+ZVx5KeIPzhcew/iBRfOjBH/dryiqAqyGKjrDjLey49hZnMD
eN4bCQNTBntZuvlpeCD9k4o8TGlVLZFE4MTyIftfQO5Vw1bMUPRodQV65AdBusnS
nJLQPDw7tIXZVQb+LsqSo0EMskXbfA4yddSsnEdin5Xy8tjFvZhhha8XnBDiQ5ln
eHOtZ47IECusBqwJdTwn2XB3sVifTimJaMi9rnCdOXOBl6jXFk+Kccf52fk+FRDx
1u36K2PuW/zUeifNm2JMaDglObb5Wpuyc7gabNqeUKdHBYNVXZ5rpVIedINC0qDH
AJbQxI2KNViW6wGDUN4UpMf8wQgH36A2tWjfm+ixE2Lfo5C/NO8jBBJ4CrCwdeMn
sW6VEVIkt0t8CeWue+XmnhXUoh72P+b/256VSaRuRAznlUzzKi660I+wf+4aVkJZ
aKr7VnSDeAG/JoxVfXN9cyVA6U5kshGbWj9W4nC7UjnlV8Vbuq0fv4th7izVgeCn
w2+k8YfwfDW4X2i0cYiCdqGB/GLiUp+dcCKgZPwNFD8PKs9oLjXLff8DoLaST5bv
P1hQMunAeJGHCUjDFfGOEaNRNy/vaiiR250xDOQ1+lbFc/0dccsm0O8Mfl+wr1gc
Bi1f0mLBh1daaHj8AaNaoaQ5jVrVpZxM9FpXlyqmC+SsFmVIYmj8UFsNCc/ZzaML
O4Y6MKrqGN6LAYN7S2sIVZWIU4HPHLRgy08jBtCAPSLW+sAtMbrp2jbO7SQC1Wjk
ahEVewwvcNWNptGldYc16SXbT04eP6cCMfx9ygChGDT90CSO7meIgGaVg2MCGba1
yeDZ0trRcF+le969lJlOTguHy5NDwG0CKUgdokeZh9EXUKMnarS0byvsSdESrV1E
+kgIosdmiebyQIxOAcmL7WkJbf2yRsl3g1ugMqAUAoFih/4h9rK4KCxNE2J9qPEQ
y/MYCzavN23f0HzDBmAtMGTKmXPtX4Zuc8nrILXgTkvb9riZFAhcJ7os/mXoUIgU
xt5i2KOlntgF6sRA53qgztFEDmhrzir4tXHEEUXWw/S8m6hzlhbmVOxYE1D5ni85
h39c+2PYSLg6ILF/sdUel1JeaLMp+4Nj5mE8iZ6Gw/WfRaGLXhbkG3RJVs5Swr8c
Og6IgjW4fKgPIoYehCKjn/9+GCSxFp/xB9gQACSHkJt9dyZTc+nCkar8TV/5S0Hz
c45tNCVYIED48RYAoj0A2Rbdz/6PZ5fUwDilzwhOozpFsDdJaEo3Ae0ErGWL2hsk
7bt1AnYu74SqxyNWqCkDbIphlfp5scZs22TRRPvzmA1eW1B1h4JU/JJCBHfEIiPq
gOQGeRH4nHGp4YJr0gSisEnCc0RH4iGkoPr1u/sflpGEiv6ZmZ+2YHdTJVARGra1
XsqPlqPZnpSsBevCyMIilfOWLkHFJLhdC4qsnGNb4TKKVx4CPqoXRMpMtbF7imXC
tiHV2pwto6Nd2wQUMy7vuZhYViOD7p6tqJ6VO2nC9In04u19KIFK/L16oMBtfN8k
kI+32KlOSqCgc2wpbC0GiHirW66Hx7klO2ygIQ0SFn2Z3VkAIXN4pcaQWycxtKLa
+aT20x4K6mcC5wYhFclrmI1UzVpyfhLXjnWGPyV6PnA0X9anXRK1qBc/d6HqSgg+
OnJDW9UgheBOS3icRfoNrTkEsAWjq9nzSuP61UZ7r7qdLUeUh8h1W15JY69JhGkv
KKawCUfVNrsuvjx/ND+SfnrU6rNRhnZysV4heV8KYRc2A5+3UugjG2vcidaLqWKP
VFdG13hmcYwlSsgZOi7syN1vj4f4KybnVjaeLfvSAlnjgO6vfi77wkfA4t6teMV9
pMOzykpkPi8o8eJQOYcOVTPEOWmmO8Eu3eV6atzj1URE/l1GzfA+MHIluyOncxw8
xl4UTo0yTNKIO88dhADX1ous2H2p5MdsrNNRpF2wv7X++P4Pj+PQVQkKYeSwKJND
KGEschneTOVwZddGttjVzwyNXrF30E2e5Qw56mx8uN1pxFyI3IzREGD/ihTmHnta
NaO4wSMaUdZobfZBwlRLwJKFiMQJ2kv4y6bLtKnFiB/mujbDt7C8NMoIdHow2vla
lDmN0ho74+s3IlzY2LVr2S4/RtYyzGtsTEojYGZsfdC9CacWFZzeqyAKSywixwFd
8ecuD8h0K2psy3zc/+TbU8pSLW78HOi+s/wmSsHA5nelt+7sNL4G59JdlOf9b90a
v6sTQLVfrBPih+xQ1L+VAC8nr5YtF4BVsLLo/ZdkjX/CoraiR+D8YLbF4zn7OXFu
Nk9QyyvyrSKiCaLER6QilwOrxaaGkThpElaxkY28KHolgH6AbLOefxb8jEEAeQWI
qksRwkFxnhBPWFYtgdErf7NQM5+U2Yr0VikrkxG2MF9CnFNw/QCfg0UlOXlK7pY7
xGgodmyWL4AgvDELWZPMNNq4tbzsfGOavg4vpYmyV61BpmhLJupJpnFhsLuLztHx
0+3BOHLzw8wa+YXPehLt8Gqa0csLiYki2KsCA00dSa47UJ2+V/8A7EzrD76R3qYo
Kr0Q9kDztA+6h9ZwiM4QcAblW8cROU1XvHmPmrzFAJG4opMF/of0uhWvIyz9V1IX
hRio6xz26VOAaj7JvATbYRLeEGhc6SeXH9EBVPDLVerbMeMV4rlC4D/Wip0eSAk0
CEhnCRK6lgnlv/7L3tPYqGiWtNTzpy+myoJHua/FJX6HX+VAVL11qzaVC3rnmEKq
zvjFldrZlCnu7uXyz9CcmlzQEXxgYOH81R8naRB7gxngfW6cBYnycYlLOpz0uFH0
z5HSFd/ym9+c7Mh+3h8UeO3r5/jAwvCrJ/tb6HHrbtBiutZG7Vp7r405ei5twVxL
7oGcfQz/GLF5H81mpnOPEfHFWWKsyQzrGyICAFrGXJT81QBiXmTCmUAV/TuxKpWu
RaIzqoqAjhq3km8d1O8T6GR672RIcm58SHNH4wEo2CBznkmlKIxL2pO+ynyw85L8
EiUSO+MgRRFLCj/edu+LHJWQiee+VWs1XwB42u6V/ZovGuxxhgnbPb4CbBp5GFuS
u3BxW2HtRi0VKPMq20WsPVb7QfWMsh5+QXzou7D0Z5SSmEiPxGY1iHMF2bAKnvJb
WBlwY5+Eg3W/8+hiB3gqintVTKSOGwGuwWpJXxuMMJE1Fgm3ZuIyckE/NBbS1DkD
XQE8IxBEArJWwyRCOPlsT2PQNu+4LJxhuNLLpNMosTfSd7tDha2TZc2MpDqJQjNY
UP6H9JUgV2LAT5YwdURL0wQa0V62TAk0WPOBSGujxkJ9gyMw2nlNhiLbkeeEfwqz
0aKzlytobS7iJphlVQcBTyWFNPYrZkfdj2WtaHLfRU3DR0s6SdWKXAy1MVB5R80p
VpHc7vPBSnNKsrPpfzpl6hF3tfeUAV0OvxF5KidTkbkfNlj+PZ2y/XXWCZ4kA05I
HFobkG17eixg7xHOn5qd01egDK9fyeDiUAgx+iWYojBbWSYpvqX0TByFNJSet3Y6
v/dTNvyX7vlJIPZ+EZJ0KWS6175zfbbd9VBdcsDow1VjzZLqlLSQO7lKsAwue06l
stxelE468NzO0d8ZkLSBf4Z61cSQVUlTsrOS1W0VLpqf0MPt3PVmUTh/wz7KZxMK
DQtrITJb7ysF2eaL6kVV5oFJtwaP7iEaKhUXHDAQQb1ezwgSdnNEUQ1Iv+Jin9SC
SnGE0Op9D5ODWkRWzU18tXcqmRK6+ZQRinRwBddrv9aZlWAApatxKfGOru2B9uFW
2bJvhfLVCguEtN2Wy+9jdcvkEoHAhY3dEN3LyjaX/7CCv0WwM26XJ7od41N809xl
NL3GryxqBUW3mlgtNkdCyGOAWXuV+y0MLUubpoAd6zCzmnYbJMs1fzafK+9UIsDY
tPkUXz2i21LVq2wWDRNfYMDz6NY5n0ncp1LzRkFpFwnnNWvZLMeGV/0LHNPcYgD2
QUiljDcjq/qx8CzVIPCXwGNHWvt88FYrZKPyl2o1inWosH4e1UMOdwrJzAP9JWfn
rynNU2j/WDzTBSMd1EnFGA5kegqdZQLRx35qf4nzSt+8puw97/yIFS8PkomkRJnz
BJdzCAymCBs4fshYx4chFCIVqL/rjrJ0RX1AFiEwryZ42e+SN5Pfs2+VedjppRUP
t4p39ewUx1hs1p4sBqa1reR5MNkPpeUatJtsQzkP95nDpR46sXEWO8yqcQJf7ECM
1QGvFnj/J+mfOwtZRzAxHcBXtTlM3AOZQirO0HxusdZphPVYKW9qPg2mmyaxXpfS
rbCN5o/PUYfMk1MM0NTfydgM6J6Ut9dWxR6rbTpwrFrPWeJYqX2TUKCaCR60UOGS
qKk46YWKK1UmeWnaOT9/nMenpXxKKx4/agGNBZw5+CDcGmJSx+rJwzrw9id2z0Fs
HFqQr06wUX/KZHneQ2t6mF1pTJNbKAah5pNZz6xZibnXW2p7bDX/2wnA/ZT5xMYR
1I3hch2ALlrUNQmpFRrbQ0PkXkgkXXzlY6uTeJN1mpkMAjZZ6gMbE3WTRUf+yIPm
ZdsDlcPgxnKA8laWAsNhPEKn6t2pzBIHdgX/A5z55L1CalYP0splo/j/aPNHzzaj
0pcx2lCyMuXdCYsIJ7rkmXwDA5Sz1iXckThoq5gJIHSlWnkFOXQvdgMBQ7cgKgE8
h6nviaQmuQstSxEo5DeTe31K+9zoQvLLm6xUv5vsw3n/MQg9TGDBuRv3+hUvhVUh
IZY21KXL7rZufLbAzw7X9/H3l3mFkYoJQXiVdT3RM0HbziQH6iCXWIIc8biOTeQb
vO/VMBgMiP/wdaL1PWHsAFobdKdH8/uEEtG9q+GYFhFPWPtTZcy7wlGTtVvjcEVF
8aDX7Ckke4accLnViyDsh6f4t8uu0ls++loV0sBQgzA0NPUDICPtCVdU+aoT3qhJ
Dgzvjpz5/79URhIzlqmXXnhCS4h7MBfu/7IfzEZh/4mCs8g7eAbqbXy+mxKdkME4
X2ck2Lkyw8cLV+6JUde7nvR9He9invilwGPzIJWANuCFgQ30gakTCGpzVJBNnb+t
v5P5bPVCdOF4kUpVDS6Mg2NhDXVJXNkVGpbAq3+IzWku7omiH++35BljFa+T91KJ
wJ7J0/P+IZ7HJx8L3+AhdnRcHxIw9C6MharTXUy2VQTDS7DR8caCGbeD6JOQGm+F
H0fq4ZlhVMNRaR2JeXfffwdtkrEo5ue4JkbztJg+iJi1T59Tse0D7TZ3ssfHX+l3
819kNyeT7rYRLjdej3NOunOLlyscHVQz75GbnAaPQ7Y9V+LVgH3+3whuWjgfY9hr
kBQgS51ZwBWHJvueeHoVovHDHrlmff7o8h9pqvJ8CZ5onUMs21r7GxuJB9JAWqin
W1ZjbIvr4aoCS7r2QIi/QReJA0WH7eHZgwL+aA1ngsLbSXPBR0Yt2A4AqMMeFef6
PfSgWfy+58exyp1w+Fu6/c1AbLv+QtfJsBovoJhLxSz9LkfRhkaqgyzt6kW+RZGk
i9NMHzZQBYyqhfLFyVqf3H/WSq9AgqIE5kwG5b/V4aghiOvPq1CV+pFVkxPwBcK9
aCfKg023fExt2fFgfgXnFWePmUuLPDzrRKKG/AA8nZExthfohltTNWKId8/OmR2d
VSXr21KtyMJmiuGmHGAnZXG5J+BfjomeLh/eGDjjthKUuJnuzBhngrasl60Go7AG
mvFCJYeKQ3aJy4olxIZw79iXudva8S0IGSjkAmbWyQdgBum9xrFfy8f+1I6FNIDn
nFZHJBzopRb2TOYL2FjkV/rLFBcIRRp5bKMRHalw8j+C3iTksWDu1GOgve+0QApI
kMdB50xBawXIzNzvTxneh6jZoaSh4Uipu3PtaMY94imwMXSqLYk/Em4wHT9YA4bv
r35kGunbhI7Snq7Y6Nj+GcLYkeCu/mtjBGe1WS4RkMe15Jssiez7k3fueHGSo97k
KHNgQsFmIdyf77gpXlE+OlInczughp/dH+UthOsaoqsSQuWlBtXZpT1Xv68ycEEh
4177rsPjwLdxrCvX9Z8bWoR6l60mvHxCcDeGxDrZkwY+xUs7iiBBTKdTkHbIvfYw
OCXHQcqMutQzr28JsFM6l9CejJt+dCp5BCmd3D5AYgC3gngNlQWdXUTjQF/6pjKv
tEpZjNSCmusNCFLpxIvorUHBZDSEH47ijMtoVux3Av6mxzPQamcQeDlPDmIHBb2k
glTKe1+7zKOPmnfl5t7llj+RGcRukWUXq4xZGf8wiJWzOvakOntMy3QU810VAljW
ZeOthzDgzL/kKwMy0C6zSIviuPHB52joiyUBpjP732PznkvSzCq/EkkNhkReoffd
rlEYhOPCE1JGZSeD1qmxXRIbiYuAXQ5166k83BB62mnYnf1WPsKeGMN2vrwgjjbQ
avrT79rR9f+n0HEZOuSAPvV3J07tcYq+sSjpPNcsIUu7mMW0M4w5YnICji+ZLy77
wjyIadYvEdAeCh2pIFA4UGFL9gb7HJPz9Q34DmxnL6Y=
`pragma protect end_protected
